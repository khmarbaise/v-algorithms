module main

import sorting

fn main() {
	println('Hello World!')
}