module main

import sorting

fn main() {
  nums := [7, 9, 35, 1, 12, 22]

  println('Hello World!')
  for idx, ie in nums {
    println('idx:$idx value:$ie')
  }

}