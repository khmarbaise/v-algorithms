module sorting

fn init() {
	println('Sorting Module!')
}

fn bubble_sort() {

}
