module sorting

fn init() {
	println('Sorting Module!')
}

fn bubble_sort<T>(unsorted[]T) []T {
 nums := unsorted.clone()
 return nums
}
