module assert_that

pub fn current<T>(unsorted[]T) []T{
  return []
}